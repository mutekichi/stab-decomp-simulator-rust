3.535533905932736198e-01,8.129419882081720845e-18
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
-2.499999999999998890e-01,2.499999999999998890e-01
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
3.535533905932736198e-01,-8.129419882081720845e-18
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
-2.499999999999998890e-01,2.499999999999998890e-01
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
-8.129419882081720845e-18,3.535533905932736198e-01
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
-2.499999999999998890e-01,-2.499999999999998890e-01
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
8.129419882081720845e-18,3.535533905932736198e-01
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
-2.499999999999998890e-01,-2.499999999999998890e-01
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00

-5.177669529663684461e-02,1.249999999999998612e-01
3.017766952966364769e-01,-1.249999999999998612e-01
-3.017766952966365324e-01,-1.249999999999998612e-01
5.177669529663678216e-02,1.249999999999998612e-01
1.249999999999998751e-01,-5.177669529663676828e-02
-1.249999999999998612e-01,3.017766952966364769e-01
1.249999999999998612e-01,3.017766952966365324e-01
-1.249999999999998612e-01,-5.177669529663685155e-02
-5.177669529663675441e-02,-1.249999999999997502e-01
-1.249999999999998335e-01,3.017766952966365324e-01
3.017766952966365324e-01,-1.249999999999998612e-01
-1.249999999999998612e-01,-5.177669529663683073e-02
-5.177669529663684461e-02,1.249999999999998612e-01
-1.249999999999999029e-01,-3.017766952966365879e-01
-3.017766952966365324e-01,-1.249999999999998612e-01
1.249999999999998057e-01,-5.177669529663677522e-02

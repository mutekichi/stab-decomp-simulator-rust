4.353579982418467712e-18,1.767766952966366434e-01
1.249999999999998890e-01,-3.749999999999994449e-01
1.767766952966365879e-01,2.340199563321044580e-17
-1.249999999999997780e-01,1.249999999999997780e-01
-1.249999999999997780e-01,1.249999999999998612e-01
-3.535533905932732313e-01,1.767766952966365879e-01
-1.249999999999998335e-01,-1.249999999999997780e-01
-1.767766952966365879e-01,2.775557561562891351e-17
1.767766952966365601e-01,-1.289152379477972153e-17
3.749999999999993339e-01,1.249999999999997502e-01
-1.120786581008785529e-17,-1.767766952966365324e-01
-1.249999999999997780e-01,-1.249999999999997502e-01
1.249999999999997363e-01,1.249999999999998196e-01
-1.767766952966365324e-01,-3.535533905932730647e-01
-1.249999999999997363e-01,1.249999999999997086e-01
2.775557561562891351e-17,-1.767766952966365324e-01

-1.821383476483178776e-01,-1.013325214724773160e-01
-1.562499999999996114e-01,1.013325214724772882e-01
-1.294417382415917472e-02,-1.714150429449547708e-01
3.879441738241580784e-01,3.124999999999987857e-02
9.374999999999961142e-02,-3.406092167691134875e-01
-2.705266952966361438e-01,2.004441738241585780e-01
-2.004441738241586890e-01,2.080266952966363381e-01
-1.379441738241588555e-01,-8.302669529663667114e-02
1.379441738241587445e-01,1.455266952966363936e-01
-2.004441738241586335e-01,2.705266952966361438e-01
-3.124999999999997224e-02,1.272208691207956099e-01
-2.080266952966363658e-01,1.638325214724772327e-01
-4.955582617584061017e-02,1.928616523516810677e-01
7.544417382415900819e-02,-2.705266952966359773e-01
-1.821383476483179609e-01,1.294417382415928575e-02
-2.052669529663683420e-02,1.294417382415917819e-02
